module Comand_dec (clk, rst, instruction, \disable , add, sub, \not , \or , \nor , \xor , nxor, \and , \nand , mul, div);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] instruction;
  input  wire [0:0] \disable ;
  output  wire [0:0] add;
  output  wire [0:0] sub;
  output  wire [0:0] \not ;
  output  wire [0:0] \or ;
  output  wire [0:0] \nor ;
  output  wire [0:0] \xor ;
  output  wire [0:0] nxor;
  output  wire [0:0] \and ;
  output  wire [0:0] \nand ;
  output  wire [0:0] mul;
  output  wire [0:0] div;

  TC_Splitter8 # (.UUID(64'd4482002304585879758 ^ UUID)) Splitter8_0 (.in(wire_26), .out0(wire_17), .out1(wire_3), .out2(wire_9), .out3(wire_11), .out4(), .out5(), .out6(), .out7());
  TC_And # (.UUID(64'd4252431844707396293 ^ UUID), .BIT_WIDTH(64'd1)) And_1 (.in0(wire_10), .in1(wire_4), .out(wire_5));
  TC_And # (.UUID(64'd4144751353222221780 ^ UUID), .BIT_WIDTH(64'd1)) And_2 (.in0(wire_6), .in1(wire_4), .out(wire_22));
  TC_And # (.UUID(64'd4133577518381962296 ^ UUID), .BIT_WIDTH(64'd1)) And_3 (.in0(wire_14), .in1(wire_4), .out(wire_25));
  TC_And # (.UUID(64'd1986947325099471790 ^ UUID), .BIT_WIDTH(64'd1)) And_4 (.in0(wire_0), .in1(wire_4), .out(wire_27));
  TC_And # (.UUID(64'd1658103694235915076 ^ UUID), .BIT_WIDTH(64'd1)) And_5 (.in0(wire_28), .in1(wire_4), .out(wire_7));
  TC_And # (.UUID(64'd2475509357815399716 ^ UUID), .BIT_WIDTH(64'd1)) And_6 (.in0(wire_13), .in1(wire_4), .out(wire_2));
  TC_And # (.UUID(64'd117348881111616919 ^ UUID), .BIT_WIDTH(64'd1)) And_7 (.in0(wire_20), .in1(wire_4), .out(wire_12));
  TC_And # (.UUID(64'd3536995208825527405 ^ UUID), .BIT_WIDTH(64'd1)) And_8 (.in0(wire_19), .in1(wire_4), .out(wire_18));
  TC_And # (.UUID(64'd1238735380101438541 ^ UUID), .BIT_WIDTH(64'd1)) And_9 (.in0(wire_21), .in1(wire_4), .out(wire_8));
  TC_And # (.UUID(64'd4146951805569167914 ^ UUID), .BIT_WIDTH(64'd1)) And_10 (.in0(wire_23), .in1(wire_4), .out(wire_1));
  TC_And # (.UUID(64'd634370225490012296 ^ UUID), .BIT_WIDTH(64'd1)) And_11 (.in0(wire_24), .in1(wire_4), .out(wire_16));
  _4bit_decoder # (.UUID(64'd1146183311277553230 ^ UUID)) _4bit_decoder_12 (.clk(clk), .rst(rst), .\1_Bit (wire_17), .\3_Bit (wire_9), .\4_Bit (wire_11), .\2_Bit (wire_3), .\16 (), .\1 (wire_10), .\2 (wire_6), .\3 (wire_14), .\4 (wire_0), .\5 (wire_28), .\7 (wire_20), .\8 (wire_19), .\9 (wire_21), .\10 (wire_23), .\11 (wire_24), .\12 (), .\13 (), .\14 (), .\15 (), .\6 (wire_13));
  TC_Not # (.UUID(64'd3630807895362982839 ^ UUID), .BIT_WIDTH(64'd1)) Not_13 (.in(wire_15), .out(wire_4));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  assign mul = wire_1;
  wire [0:0] wire_2;
  assign \xor  = wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  assign add = wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  assign \nor  = wire_7;
  wire [0:0] wire_8;
  assign \nand  = wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  assign nxor = wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  assign wire_15 = \disable ;
  wire [0:0] wire_16;
  assign div = wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  assign \and  = wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  assign sub = wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  assign \not  = wire_25;
  wire [7:0] wire_26;
  assign wire_26 = instruction;
  wire [0:0] wire_27;
  assign \or  = wire_27;
  wire [0:0] wire_28;

endmodule
