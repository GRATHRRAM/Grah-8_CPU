module grahzm8 (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_Program # (.UUID(64'd3141827013512232805 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_2B9A0305CE1F7F65.w8.bin"), .ARG_SIG("Program_2B9A0305CE1F7F65=%s")) Program_0 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_36 }), .out0(wire_6), .out1(), .out2(), .out3());
  TC_Ram # (.UUID(64'd1442474303503021395 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_1 (.clk(clk), .rst(rst), .load(wire_34), .save(wire_3), .address({{24{1'b0}}, wire_5 }), .in0(wire_4), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_4_0), .out1(), .out2(), .out3());
  TC_Counter # (.UUID(64'd932762492408994202 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_2 (.clk(clk), .rst(rst), .save(wire_45), .in(wire_4[7:0]), .out(wire_36));
  TC_Switch # (.UUID(64'd3960965275402640681 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_3 (.en(wire_7), .in(wire_6[7:0]), .out(wire_4_8[7:0]));
  TC_Splitter8 # (.UUID(64'd1794847357655579608 ^ UUID)) Splitter8_4 (.in(wire_6[7:0]), .out0(wire_17), .out1(wire_31), .out2(wire_0), .out3(wire_13), .out4(wire_1), .out5(wire_41), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd4611564000427626573 ^ UUID)) Decoder3_5 (.dis(wire_22), .sel0(wire_13), .sel1(wire_1), .sel2(wire_41), .out0(wire_44), .out1(wire_32), .out2(wire_38), .out3(wire_26), .out4(wire_14), .out5(wire_35), .out6(wire_34), .out7(wire_28));
  TC_Decoder3 # (.UUID(64'd3975716302527489394 ^ UUID)) Decoder3_6 (.dis(wire_22), .sel0(wire_17), .sel1(wire_31), .sel2(wire_0), .out0(wire_27), .out1(wire_12), .out2(wire_16), .out3(wire_42), .out4(wire_8), .out5(wire_20), .out6(wire_3), .out7(wire_39));
  TC_Not # (.UUID(64'd2085913829163953837 ^ UUID), .BIT_WIDTH(64'd1)) Not_7 (.in(wire_37), .out(wire_22));
  TC_Switch # (.UUID(64'd592641017123523600 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_8 (.en(wire_10), .in(wire_24), .out(wire_4_4[7:0]));
  TC_Or # (.UUID(64'd2664153464624268752 ^ UUID), .BIT_WIDTH(64'd1)) Or_9 (.in0(wire_42), .in1(wire_10), .out(wire_30));
  TC_Switch # (.UUID(64'd2384141649022815990 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_10 (.en(wire_28), .in({{7{1'b0}}, wire_9 }), .out(wire_4_2[7:0]));
  TC_Switch # (.UUID(64'd1881273207972279230 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_39), .in(wire_4[7:0]), .out(wire_2));
  TC_Decoder1 # (.UUID(64'd1204120349862430746 ^ UUID)) Decoder1_12 (.sel(wire_17), .out0(wire_18), .out1(wire_25));
  TC_And # (.UUID(64'd4109806387476150794 ^ UUID), .BIT_WIDTH(64'd1)) And_13 (.in0(wire_19), .in1(wire_18), .out(wire_33));
  TC_And # (.UUID(64'd676486280697974606 ^ UUID), .BIT_WIDTH(64'd1)) And_14 (.in0(wire_25), .in1(wire_19), .out(wire_23));
  TC_Or # (.UUID(64'd1756542076950970648 ^ UUID), .BIT_WIDTH(64'd1)) Or_15 (.in0(wire_7), .in1(wire_27), .out(wire_21));
  TC_Or # (.UUID(64'd2242600398968762306 ^ UUID), .BIT_WIDTH(64'd1)) Or_16 (.in0(wire_33), .in1(wire_44), .out(wire_15));
  TC_Or # (.UUID(64'd950621913437045215 ^ UUID), .BIT_WIDTH(64'd1)) Or_17 (.in0(wire_23), .in1(wire_35), .out(wire_29));
  TC_Or # (.UUID(64'd3542487319000578313 ^ UUID), .BIT_WIDTH(64'd1)) Or_18 (.in0(wire_23), .in1(wire_33), .out(wire_45));
  TC_Switch # (.UUID(64'd1621303180505943999 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_10), .in(wire_6[7:0]), .out(wire_40));
  RegisterPlus # (.UUID(64'd2515007776148876636 ^ UUID)) RegisterPlus_20 (.clk(clk), .rst(rst), .Load(wire_15), .Save_value(wire_4[7:0]), .Save(wire_21), .Always_output(), .Output(wire_4_9[7:0]));
  RegisterPlus # (.UUID(64'd1145908529650350723 ^ UUID)) RegisterPlus_21 (.clk(clk), .rst(rst), .Load(wire_32), .Save_value(wire_4[7:0]), .Save(wire_12), .Always_output(wire_11), .Output(wire_4_7[7:0]));
  RegisterPlus # (.UUID(64'd289786154161998413 ^ UUID)) RegisterPlus_22 (.clk(clk), .rst(rst), .Load(wire_38), .Save_value(wire_4[7:0]), .Save(wire_16), .Always_output(wire_43), .Output(wire_4_6[7:0]));
  RegisterPlus # (.UUID(64'd1917400086359645051 ^ UUID)) RegisterPlus_23 (.clk(clk), .rst(rst), .Load(wire_26), .Save_value(wire_4[7:0]), .Save(wire_30), .Always_output(), .Output(wire_4_5[7:0]));
  Instruction_dec # (.UUID(64'd4582718711987810921 ^ UUID)) Instruction_dec_24 (.clk(clk), .rst(rst), .Input(wire_6[7:0]), .Val_2_Reg0(wire_7), .Copy(wire_37), .Calculate(wire_10), .Counter_Man(wire_19));
  Grahzm8_Alu # (.UUID(64'd2732743794862348741 ^ UUID)) Grahzm8_Alu_25 (.clk(clk), .rst(rst), .Input_1(wire_11), .Input_2(wire_43), .Instruction(wire_40), .Output(wire_24));
  RegisterPlus # (.UUID(64'd2399782736842396036 ^ UUID)) RegisterPlus_26 (.clk(clk), .rst(rst), .Load(wire_14), .Save_value(wire_4[7:0]), .Save(wire_8), .Always_output(wire_5), .Output(wire_4_3[7:0]));
  RegisterPlus # (.UUID(64'd4127468653178353900 ^ UUID)) RegisterPlus_27 (.clk(clk), .rst(rst), .Load(wire_29), .Save_value(wire_4[7:0]), .Save(wire_20), .Always_output(), .Output(wire_4_1[7:0]));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [7:0] wire_2;
  wire [0:0] wire_3;
  wire [63:0] wire_4;
  wire [63:0] wire_4_0;
  wire [63:0] wire_4_1;
  wire [63:0] wire_4_2;
  wire [63:0] wire_4_3;
  wire [63:0] wire_4_4;
  wire [63:0] wire_4_5;
  wire [63:0] wire_4_6;
  wire [63:0] wire_4_7;
  wire [63:0] wire_4_8;
  wire [63:0] wire_4_9;
  assign wire_4 = wire_4_0|wire_4_1|wire_4_2|wire_4_3|wire_4_4|wire_4_5|wire_4_6|wire_4_7|wire_4_8|wire_4_9;
  wire [7:0] wire_5;
  wire [63:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  assign wire_9 = 0;
  wire [0:0] wire_10;
  wire [7:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [7:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [7:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [7:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [7:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;

endmodule
