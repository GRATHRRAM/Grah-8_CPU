module _4bit_decoder (clk, rst, \1_Bit , \3_Bit , \4_Bit , \2_Bit , \16 , \1 , \2 , \3 , \4 , \5 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \6 );
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] \1_Bit ;
  input  wire [0:0] \3_Bit ;
  input  wire [0:0] \4_Bit ;
  input  wire [0:0] \2_Bit ;
  output  wire [0:0] \16 ;
  output  wire [0:0] \1 ;
  output  wire [0:0] \2 ;
  output  wire [0:0] \3 ;
  output  wire [0:0] \4 ;
  output  wire [0:0] \5 ;
  output  wire [0:0] \7 ;
  output  wire [0:0] \8 ;
  output  wire [0:0] \9 ;
  output  wire [0:0] \10 ;
  output  wire [0:0] \11 ;
  output  wire [0:0] \12 ;
  output  wire [0:0] \13 ;
  output  wire [0:0] \14 ;
  output  wire [0:0] \15 ;
  output  wire [0:0] \6 ;

  TC_Not # (.UUID(64'd4022553707154021137 ^ UUID), .BIT_WIDTH(64'd1)) Not_0 (.in(wire_6), .out(wire_32));
  TC_Not # (.UUID(64'd2504430404737194098 ^ UUID), .BIT_WIDTH(64'd1)) Not_1 (.in(wire_0), .out(wire_46));
  TC_Not # (.UUID(64'd2981285277316280103 ^ UUID), .BIT_WIDTH(64'd1)) Not_2 (.in(wire_1), .out(wire_11));
  TC_Not # (.UUID(64'd883831078267320792 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_5), .out(wire_13));
  TC_Not # (.UUID(64'd1807726004133460370 ^ UUID), .BIT_WIDTH(64'd1)) Not_4 (.in(wire_0), .out(wire_21));
  TC_Not # (.UUID(64'd1447287332920659867 ^ UUID), .BIT_WIDTH(64'd1)) Not_5 (.in(wire_1), .out(wire_2));
  TC_Not # (.UUID(64'd3161590505079411770 ^ UUID), .BIT_WIDTH(64'd1)) Not_6 (.in(wire_5), .out(wire_14));
  TC_Not # (.UUID(64'd2088207711814206694 ^ UUID), .BIT_WIDTH(64'd1)) Not_7 (.in(wire_1), .out(wire_42));
  TC_Not # (.UUID(64'd983467647963475849 ^ UUID), .BIT_WIDTH(64'd1)) Not_8 (.in(wire_5), .out(wire_4));
  TC_Not # (.UUID(64'd845581792190483065 ^ UUID), .BIT_WIDTH(64'd1)) Not_9 (.in(wire_1), .out(wire_35));
  TC_Not # (.UUID(64'd792929086023444613 ^ UUID), .BIT_WIDTH(64'd1)) Not_10 (.in(wire_5), .out(wire_3));
  TC_Not # (.UUID(64'd2451376733646595199 ^ UUID), .BIT_WIDTH(64'd1)) Not_11 (.in(wire_0), .out(wire_41));
  TC_Not # (.UUID(64'd2651844577442475059 ^ UUID), .BIT_WIDTH(64'd1)) Not_12 (.in(wire_5), .out(wire_10));
  TC_Not # (.UUID(64'd2810718856234171282 ^ UUID), .BIT_WIDTH(64'd1)) Not_13 (.in(wire_0), .out(wire_45));
  TC_Not # (.UUID(64'd2363532353380720241 ^ UUID), .BIT_WIDTH(64'd1)) Not_14 (.in(wire_5), .out(wire_44));
  TC_Not # (.UUID(64'd3415245668154633256 ^ UUID), .BIT_WIDTH(64'd1)) Not_15 (.in(wire_5), .out(wire_23));
  TC_Not # (.UUID(64'd3997128288643024462 ^ UUID), .BIT_WIDTH(64'd1)) Not_16 (.in(wire_5), .out(wire_36));
  TC_Not # (.UUID(64'd723066936421833634 ^ UUID), .BIT_WIDTH(64'd1)) Not_17 (.in(wire_0), .out(wire_48));
  TC_Not # (.UUID(64'd2137048554743263637 ^ UUID), .BIT_WIDTH(64'd1)) Not_18 (.in(wire_1), .out(wire_34));
  TC_Not # (.UUID(64'd2080220701292213205 ^ UUID), .BIT_WIDTH(64'd1)) Not_19 (.in(wire_0), .out(wire_9));
  TC_Not # (.UUID(64'd984152951232000238 ^ UUID), .BIT_WIDTH(64'd1)) Not_20 (.in(wire_1), .out(wire_18));
  TC_Not # (.UUID(64'd3339112747147205643 ^ UUID), .BIT_WIDTH(64'd1)) Not_21 (.in(wire_1), .out(wire_22));
  TC_Not # (.UUID(64'd2954264011593770418 ^ UUID), .BIT_WIDTH(64'd1)) Not_22 (.in(wire_1), .out(wire_20));
  TC_Not # (.UUID(64'd1261308213207646075 ^ UUID), .BIT_WIDTH(64'd1)) Not_23 (.in(wire_0), .out(wire_25));
  TC_Not # (.UUID(64'd1309824771915995550 ^ UUID), .BIT_WIDTH(64'd1)) Not_24 (.in(wire_0), .out(wire_51));
  TC_Not # (.UUID(64'd2445136097262996103 ^ UUID), .BIT_WIDTH(64'd1)) Not_25 (.in(wire_6), .out(wire_31));
  TC_Not # (.UUID(64'd103577521702413013 ^ UUID), .BIT_WIDTH(64'd1)) Not_26 (.in(wire_6), .out(wire_19));
  TC_Not # (.UUID(64'd508999947213099209 ^ UUID), .BIT_WIDTH(64'd1)) Not_27 (.in(wire_6), .out(wire_39));
  TC_Not # (.UUID(64'd1791580953363036799 ^ UUID), .BIT_WIDTH(64'd1)) Not_28 (.in(wire_6), .out(wire_29));
  TC_Not # (.UUID(64'd3645001039097645942 ^ UUID), .BIT_WIDTH(64'd1)) Not_29 (.in(wire_6), .out(wire_30));
  TC_Not # (.UUID(64'd4399270207851746718 ^ UUID), .BIT_WIDTH(64'd1)) Not_30 (.in(wire_6), .out(wire_8));
  TC_Not # (.UUID(64'd3480327844175439948 ^ UUID), .BIT_WIDTH(64'd1)) Not_31 (.in(wire_6), .out(wire_47));
  _4InAnd # (.UUID(64'd1881669726319765518 ^ UUID)) _4InAnd_32 (.clk(clk), .rst(rst), .Input_1(wire_32), .Input_2(wire_11), .Input_3(wire_13), .Input_4(wire_46), .Output(wire_26));
  _4InAnd # (.UUID(64'd3154201268365375329 ^ UUID)) _4InAnd_33 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_2), .Input_3(wire_14), .Input_4(wire_21), .Output(wire_16));
  _4InAnd # (.UUID(64'd682568861334433799 ^ UUID)) _4InAnd_34 (.clk(clk), .rst(rst), .Input_1(wire_31), .Input_2(wire_42), .Input_3(wire_4), .Input_4(wire_0), .Output(wire_37));
  _4InAnd # (.UUID(64'd603078280254923757 ^ UUID)) _4InAnd_35 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_35), .Input_3(wire_3), .Input_4(wire_0), .Output(wire_40));
  _4InAnd # (.UUID(64'd1008559417439783936 ^ UUID)) _4InAnd_36 (.clk(clk), .rst(rst), .Input_1(wire_19), .Input_2(wire_1), .Input_3(wire_10), .Input_4(wire_41), .Output(wire_43));
  _4InAnd # (.UUID(64'd4160003391264076492 ^ UUID)) _4InAnd_37 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_1), .Input_3(wire_44), .Input_4(wire_45), .Output(wire_33));
  _4InAnd # (.UUID(64'd3864627739082115735 ^ UUID)) _4InAnd_38 (.clk(clk), .rst(rst), .Input_1(wire_39), .Input_2(wire_1), .Input_3(wire_23), .Input_4(wire_0), .Output(wire_17));
  _4InAnd # (.UUID(64'd2030081743972221641 ^ UUID)) _4InAnd_39 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_1), .Input_3(wire_36), .Input_4(wire_0), .Output(wire_12));
  _4InAnd # (.UUID(64'd582214723974831901 ^ UUID)) _4InAnd_40 (.clk(clk), .rst(rst), .Input_1(wire_29), .Input_2(wire_34), .Input_3(wire_5), .Input_4(wire_48), .Output(wire_49));
  _4InAnd # (.UUID(64'd1580426462405451430 ^ UUID)) _4InAnd_41 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_18), .Input_3(wire_5), .Input_4(wire_9), .Output(wire_28));
  _4InAnd # (.UUID(64'd3490086501885240065 ^ UUID)) _4InAnd_42 (.clk(clk), .rst(rst), .Input_1(wire_30), .Input_2(wire_22), .Input_3(wire_5), .Input_4(wire_0), .Output(wire_24));
  _4InAnd # (.UUID(64'd774261423034419192 ^ UUID)) _4InAnd_43 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_20), .Input_3(wire_5), .Input_4(wire_0), .Output(wire_50));
  _4InAnd # (.UUID(64'd2163010496997179678 ^ UUID)) _4InAnd_44 (.clk(clk), .rst(rst), .Input_1(wire_8), .Input_2(wire_1), .Input_3(wire_5), .Input_4(wire_25), .Output(wire_7));
  _4InAnd # (.UUID(64'd4057707661934331460 ^ UUID)) _4InAnd_45 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_1), .Input_3(wire_5), .Input_4(wire_51), .Output(wire_15));
  _4InAnd # (.UUID(64'd3637058070027206394 ^ UUID)) _4InAnd_46 (.clk(clk), .rst(rst), .Input_1(wire_47), .Input_2(wire_1), .Input_3(wire_5), .Input_4(wire_0), .Output(wire_38));
  _4InAnd # (.UUID(64'd2312131805332501143 ^ UUID)) _4InAnd_47 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_1), .Input_3(wire_5), .Input_4(wire_0), .Output(wire_27));

  wire [0:0] wire_0;
  assign wire_0 = \2_Bit ;
  wire [0:0] wire_1;
  assign wire_1 = \3_Bit ;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  assign wire_5 = \4_Bit ;
  wire [0:0] wire_6;
  assign wire_6 = \1_Bit ;
  wire [0:0] wire_7;
  assign \13  = wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  assign \8  = wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  assign \14  = wire_15;
  wire [0:0] wire_16;
  assign \2  = wire_16;
  wire [0:0] wire_17;
  assign \7  = wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  assign \11  = wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  assign \1  = wire_26;
  wire [0:0] wire_27;
  assign \16  = wire_27;
  wire [0:0] wire_28;
  assign \10  = wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  assign \6  = wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  assign \3  = wire_37;
  wire [0:0] wire_38;
  assign \15  = wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  assign \4  = wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  assign \5  = wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  assign \9  = wire_49;
  wire [0:0] wire_50;
  assign \12  = wire_50;
  wire [0:0] wire_51;

endmodule
